//Add verif code here
