//Add code for corresponding code
interface  uvm_test_if;
  
endinterface
