//Add code for corresponding code
interface  uvm_test_if;
  bit[7:0] input_a;
  bit[7:0] input_b;
  bit      input_sel;
  bit[7:0] output_y
  
endinterface
