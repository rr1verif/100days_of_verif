//Agent file is used to create instance of monitor, driver and sequencer (if active agent then driver and sequencer is created")
