package uvm_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.sv"
  //Add any define file required `include 
  `include "uvm_env.sv"
endpackage
